VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO SRAM_32x128_1rw
   CLASS BLOCK ;
   SIZE 138.11 BY 75.235 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.8425 0.0 30.9825 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.7025 0.0 33.8425 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.5625 0.0 36.7025 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.4225 0.0 39.5625 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.2825 0.0 42.4225 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.1425 0.0 45.2825 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.0025 0.0 48.1425 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.8625 0.0 51.0025 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.7225 0.0 53.8625 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.5825 0.0 56.7225 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.4425 0.0 59.5825 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.3025 0.0 62.4425 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.1625 0.0 65.3025 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.0225 0.0 68.1625 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.8825 0.0 71.0225 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.7425 0.0 73.8825 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.6025 0.0 76.7425 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.4625 0.0 79.6025 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.3225 0.0 82.4625 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.1825 0.0 85.3225 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.0425 0.0 88.1825 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.9025 0.0 91.0425 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.7625 0.0 93.9025 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.6225 0.0 96.7625 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.4825 0.0 99.6225 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.3425 0.0 102.4825 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  105.2025 0.0 105.3425 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.0625 0.0 108.2025 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.9225 0.0 111.0625 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.7825 0.0 113.9225 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.6425 0.0 116.7825 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.5025 0.0 119.6425 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  25.1225 0.0 25.2625 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.9825 0.0 28.1225 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 46.99 0.14 47.13 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 49.72 0.14 49.86 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 51.93 0.14 52.07 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 54.66 0.14 54.8 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  19.405 75.095 19.545 75.235 ;
      END
   END addr0[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 5.0 0.14 5.14 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 7.73 0.14 7.87 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.84 0.0 9.98 0.14 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.9125 0.0 43.0525 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.7325 0.0 45.8725 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  48.5525 0.0 48.6925 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.3725 0.0 51.5125 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.1925 0.0 54.3325 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  57.0125 0.0 57.1525 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.8325 0.0 59.9725 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.6525 0.0 62.7925 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.4725 0.0 65.6125 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.3075 0.0 68.4475 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  71.185 0.0 71.325 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  74.0275 0.0 74.1675 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.8875 0.0 77.0275 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.7475 0.0 79.8875 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.6075 0.0 82.7475 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.4675 0.0 85.6075 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  88.3275 0.0 88.4675 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  91.1875 0.0 91.3275 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  94.245 0.0 94.385 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  97.065 0.0 97.205 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.885 0.0 100.025 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.585 0.0 101.725 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.445 0.0 104.585 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.305 0.0 107.445 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.165 0.0 110.305 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.025 0.0 113.165 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  115.885 0.0 116.025 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  118.745 0.0 118.885 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  121.605 0.0 121.745 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  124.6925 0.0 124.8325 0.14 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.97 13.1625 138.11 13.3025 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  137.97 12.9275 138.11 13.0675 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 138.11 0.7 ;
         LAYER metal4 ;
         RECT  137.41 0.0 138.11 75.235 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 75.235 ;
         LAYER metal3 ;
         RECT  0.0 74.535 138.11 75.235 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.4 1.4 136.71 2.1 ;
         LAYER metal3 ;
         RECT  1.4 73.135 136.71 73.835 ;
         LAYER metal4 ;
         RECT  136.01 1.4 136.71 73.835 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 73.835 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 137.97 75.095 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 137.97 75.095 ;
   LAYER  metal3 ;
      RECT  0.28 46.85 137.97 47.27 ;
      RECT  0.14 47.27 0.28 49.58 ;
      RECT  0.14 50.0 0.28 51.79 ;
      RECT  0.14 52.21 0.28 54.52 ;
      RECT  0.14 5.28 0.28 7.59 ;
      RECT  0.14 8.01 0.28 46.85 ;
      RECT  0.28 13.0225 137.83 13.4425 ;
      RECT  0.28 13.4425 137.83 46.85 ;
      RECT  137.83 13.4425 137.97 46.85 ;
      RECT  0.14 0.84 0.28 4.86 ;
      RECT  137.83 0.84 137.97 12.7875 ;
      RECT  0.14 54.94 0.28 74.395 ;
      RECT  0.28 0.84 1.26 1.26 ;
      RECT  0.28 1.26 1.26 2.24 ;
      RECT  0.28 2.24 1.26 13.0225 ;
      RECT  1.26 0.84 136.85 1.26 ;
      RECT  1.26 2.24 136.85 13.0225 ;
      RECT  136.85 0.84 137.83 1.26 ;
      RECT  136.85 1.26 137.83 2.24 ;
      RECT  136.85 2.24 137.83 13.0225 ;
      RECT  0.28 47.27 1.26 72.995 ;
      RECT  0.28 72.995 1.26 73.975 ;
      RECT  0.28 73.975 1.26 74.395 ;
      RECT  1.26 47.27 136.85 72.995 ;
      RECT  1.26 73.975 136.85 74.395 ;
      RECT  136.85 47.27 137.97 72.995 ;
      RECT  136.85 72.995 137.97 73.975 ;
      RECT  136.85 73.975 137.97 74.395 ;
   LAYER  metal4 ;
      RECT  30.5625 0.42 31.2625 75.095 ;
      RECT  31.2625 0.14 33.4225 0.42 ;
      RECT  34.1225 0.14 36.2825 0.42 ;
      RECT  36.9825 0.14 39.1425 0.42 ;
      RECT  39.8425 0.14 42.0025 0.42 ;
      RECT  25.5425 0.14 27.7025 0.42 ;
      RECT  28.4025 0.14 30.5625 0.42 ;
      RECT  19.125 0.42 19.825 74.815 ;
      RECT  19.825 0.42 30.5625 74.815 ;
      RECT  19.825 74.815 30.5625 75.095 ;
      RECT  10.26 0.14 24.8425 0.42 ;
      RECT  43.3325 0.14 44.8625 0.42 ;
      RECT  46.1525 0.14 47.7225 0.42 ;
      RECT  48.9725 0.14 50.5825 0.42 ;
      RECT  51.7925 0.14 53.4425 0.42 ;
      RECT  54.6125 0.14 56.3025 0.42 ;
      RECT  57.4325 0.14 59.1625 0.42 ;
      RECT  60.2525 0.14 62.0225 0.42 ;
      RECT  63.0725 0.14 64.8825 0.42 ;
      RECT  65.8925 0.14 67.7425 0.42 ;
      RECT  68.7275 0.14 70.6025 0.42 ;
      RECT  71.605 0.14 73.4625 0.42 ;
      RECT  74.4475 0.14 76.3225 0.42 ;
      RECT  77.3075 0.14 79.1825 0.42 ;
      RECT  80.1675 0.14 82.0425 0.42 ;
      RECT  83.0275 0.14 84.9025 0.42 ;
      RECT  85.8875 0.14 87.7625 0.42 ;
      RECT  88.7475 0.14 90.6225 0.42 ;
      RECT  91.6075 0.14 93.4825 0.42 ;
      RECT  94.665 0.14 96.3425 0.42 ;
      RECT  97.485 0.14 99.2025 0.42 ;
      RECT  100.305 0.14 101.305 0.42 ;
      RECT  102.005 0.14 102.0625 0.42 ;
      RECT  102.7625 0.14 104.165 0.42 ;
      RECT  104.865 0.14 104.9225 0.42 ;
      RECT  105.6225 0.14 107.025 0.42 ;
      RECT  107.725 0.14 107.7825 0.42 ;
      RECT  108.4825 0.14 109.885 0.42 ;
      RECT  110.585 0.14 110.6425 0.42 ;
      RECT  111.3425 0.14 112.745 0.42 ;
      RECT  113.445 0.14 113.5025 0.42 ;
      RECT  114.2025 0.14 115.605 0.42 ;
      RECT  116.305 0.14 116.3625 0.42 ;
      RECT  117.0625 0.14 118.465 0.42 ;
      RECT  119.165 0.14 119.2225 0.42 ;
      RECT  119.9225 0.14 121.325 0.42 ;
      RECT  122.025 0.14 124.4125 0.42 ;
      RECT  125.1125 0.14 137.13 0.42 ;
      RECT  0.98 74.815 19.125 75.095 ;
      RECT  0.98 0.14 9.56 0.42 ;
      RECT  31.2625 0.42 135.73 1.12 ;
      RECT  31.2625 1.12 135.73 74.115 ;
      RECT  31.2625 74.115 135.73 75.095 ;
      RECT  135.73 0.42 136.99 1.12 ;
      RECT  135.73 74.115 136.99 75.095 ;
      RECT  136.99 0.42 137.13 1.12 ;
      RECT  136.99 1.12 137.13 74.115 ;
      RECT  136.99 74.115 137.13 75.095 ;
      RECT  0.98 0.42 1.12 1.12 ;
      RECT  0.98 1.12 1.12 74.115 ;
      RECT  0.98 74.115 1.12 74.815 ;
      RECT  1.12 0.42 2.38 1.12 ;
      RECT  1.12 74.115 2.38 74.815 ;
      RECT  2.38 0.42 19.125 1.12 ;
      RECT  2.38 1.12 19.125 74.115 ;
      RECT  2.38 74.115 19.125 74.815 ;
   END
END    SRAM_32x128_1rw
END    LIBRARY
